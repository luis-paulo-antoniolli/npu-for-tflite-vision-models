module tflite_softcore (
    input clk,
    input rst_n,
    
    // Interface de memória unificada (multiplexada)
    input [31:0] mem_addr,
    input [31:0] mem_data_in,
    input mem_we,
    input mem_re,
    input mem_ready,
    output [31:0] mem_data_out,
    output mem_req,
    
    // Interface com NPU
    // Removed undriven signals to fix synthesis warnings
    input npu_cmd_ready,
    input [31:0] npu_result,
    input npu_result_valid,
    
    // Interface PCIe
    input [31:0] pcie_rx_data,
    input pcie_rx_valid,
    input pcie_tx_ready,
    output [31:0] pcie_tx_data,
    output pcie_tx_valid,
    
    // Sinais de status
    output [31:0] status_data,
    output [3:0] status_sel  // 0000=pc, 0001=alu_result, 0010=ready, 0011=done
);

    // Sinais de controle da NPU
    reg [31:0] npu_instruction;
    reg npu_start;
    wire npu_busy;
    
    // Pipeline de 5 estágios para melhor utilização dos recursos
    localparam FETCH = 3'b000;
    localparam DECODE = 3'b001;
    localparam EXECUTE = 3'b010;
    localparam MEMORY = 3'b011;
    localparam WRITEBACK = 3'b100;
    
    // Registradores de pipeline
    reg [31:0] pc_reg;
    reg [31:0] pc_next;
    reg [31:0] instruction_f;  // FETCH
    reg [31:0] instruction_d;  // DECODE
    reg [31:0] rs1_data_d, rs2_data_d;
    reg [4:0] rd_addr_d;
    reg [31:0] alu_a_d, alu_b_d;
    reg [3:0] alu_op_d;
    reg [1:0] imm_sel_d;
    reg pc_sel_d;
    reg alu_a_sel_d, alu_b_sel_d;
    reg mem_we_d;
    reg [1:0] wb_sel_d;
    
    reg [31:0] alu_result_e;   // EXECUTE
    reg [31:0] rs2_data_e;
    reg [4:0] rd_addr_e;
    reg mem_we_e;
    reg [1:0] wb_sel_e;
    reg zero_flag_e;
    
    reg [31:0] mem_read_data_m; // MEMORY
    reg [31:0] alu_result_m;
    reg [4:0] rd_addr_m;
    reg [1:0] wb_sel_m;
    
    reg [31:0] writeback_data_w; // WRITEBACK
    reg [4:0] rd_addr_w;
    
    // Definição dos sinais de controle
    wire [3:0] alu_op;
    wire [1:0] imm_sel;
    wire pc_sel;
    wire alu_a_sel;
    wire alu_b_sel;
    wire mem_we_ctrl;
    wire [1:0] wb_sel;
    
    // Definição dos sinais de dados
    wire [31:0] immediate;
    wire [31:0] rs1_data;
    wire [31:0] rs2_data;
    wire [31:0] alu_a;
    wire [31:0] alu_b;
    wire [31:0] alu_out;
    wire zero_flag;
    
    // Definição dos sinais de registradores
    wire [4:0] rd_addr;
    wire [4:0] rs1_addr;
    wire [4:0] rs2_addr;
    
    // Banco de registradores com dual-port read
    reg [31:0] registers [0:31];
    integer i;
    
    // Inicialização do banco de registradores
    always @(posedge clk) begin
        if (!rst_n) begin
            for (i = 0; i < 32; i = i + 1) begin
                registers[i] <= 32'h00000000;
            end
        end
    end
    
    // Pipeline: FETCH
    always @(posedge clk) begin
        if (!rst_n) begin
            pc_reg <= 32'h00000000;
            instruction_f <= 32'h00000000;
        end else begin
            pc_reg <= pc_next;
            instruction_f <= mem_data_out; // Instrução lida da memória
        end
    end
    
    // Pipeline: DECODE
    always @(posedge clk) begin
        if (!rst_n) begin
            instruction_d <= 32'h00000000;
            rs1_data_d <= 32'h00000000;
            rs2_data_d <= 32'h00000000;
            rd_addr_d <= 5'h0;
            alu_a_d <= 32'h00000000;
            alu_b_d <= 32'h00000000;
            alu_op_d <= 4'h0;
            imm_sel_d <= 2'h0;
            pc_sel_d <= 1'b0;
            alu_a_sel_d <= 1'b0;
            alu_b_sel_d <= 1'b0;
            mem_we_d <= 1'b0;
            wb_sel_d <= 2'h0;
        end else begin
            instruction_d <= instruction_f;
            rs1_data_d <= registers[instruction_f[19:15]];
            rs2_data_d <= registers[instruction_f[24:20]];
            rd_addr_d <= instruction_f[11:7];
            alu_a_d <= alu_a;
            alu_b_d <= alu_b;
            alu_op_d <= alu_op;
            imm_sel_d <= imm_sel;
            pc_sel_d <= pc_sel;
            alu_a_sel_d <= alu_a_sel;
            alu_b_sel_d <= alu_b_sel;
            mem_we_d <= mem_we_ctrl;
            wb_sel_d <= wb_sel;
        end
    end
    
    // Pipeline: EXECUTE
    always @(posedge clk) begin
        if (!rst_n) begin
            alu_result_e <= 32'h00000000;
            rs2_data_e <= 32'h00000000;
            rd_addr_e <= 5'h0;
            mem_we_e <= 1'b0;
            wb_sel_e <= 2'h0;
            zero_flag_e <= 1'b0;
            npu_start <= 1'b0;
        end else begin
            alu_result_e <= alu_out;
            rs2_data_e <= rs2_data_d;
            rd_addr_e <= rd_addr_d;
            mem_we_e <= mem_we_d;
            wb_sel_e <= wb_sel_d;
            zero_flag_e <= zero_flag;
            
            // Controle da NPU
            if (alu_op_d == 4'b1111) begin // CUSTOM instruction
                npu_start <= 1'b1;
                npu_instruction <= instruction_d;
            end else begin
                npu_start <= 1'b0;
            end
        end
    end
    
    // Pipeline: MEMORY
    always @(posedge clk) begin
        if (!rst_n) begin
            mem_read_data_m <= 32'h00000000;
            alu_result_m <= 32'h00000000;
            rd_addr_m <= 5'h0;
            wb_sel_m <= 2'h0;
        end else begin
            mem_read_data_m <= mem_data_out;
            alu_result_m <= alu_result_e;
            rd_addr_m <= rd_addr_e;
            wb_sel_m <= wb_sel_e;
        end
    end
    
    // Pipeline: WRITEBACK
    always @(posedge clk) begin
        if (!rst_n) begin
            writeback_data_w <= 32'h00000000;
            rd_addr_w <= 5'h0;
        end else begin
            writeback_data_w <= (wb_sel_m == 2'b00) ? alu_result_m :
                              (wb_sel_m == 2'b01) ? mem_read_data_m :
                              (wb_sel_m == 2'b10) ? pc_next :
                              32'h00000000;
            rd_addr_w <= rd_addr_m;
        end
    end
    
    // Escrita no banco de registradores
    always @(posedge clk) begin
        if (rd_addr_w != 5'h0) begin
            registers[rd_addr_w] <= writeback_data_w;
        end
    end
    
    // Unidade de controle
    control_unit cu (
        .opcode(instruction_d[6:0]),
        .funct3(instruction_d[14:12]),
        .funct7(instruction_d[31:25]),
        .alu_op(alu_op),
        .imm_sel(imm_sel),
        .pc_sel(pc_sel),
        .reg_we(),
        .alu_a_sel(alu_a_sel),
        .alu_b_sel(alu_b_sel),
        .mem_we(mem_we_ctrl),
        .wb_sel(wb_sel)
    );
    
    // Gerador de imediatos
    immediate_generator ig (
        .instruction(instruction_d),
        .imm_sel(imm_sel_d),
        .immediate(immediate)
    );
    
    // Seleção das entradas da ALU
    assign alu_a = alu_a_sel_d ? pc_reg : rs1_data_d;
    assign alu_b = alu_b_sel_d ? immediate : rs2_data_d;
    
    // Unidade lógica aritmética
    alu alu_inst (
        .a(alu_a_d),
        .b(alu_b_d),
        .op(alu_op_d),
        .result(alu_out),
        .zero(zero_flag)
    );
    
    // Lógica de próximo PC
    always @(*) begin
        if (pc_sel_d) begin
            // JAL
            pc_next = pc_reg + 32'h00000004;
        end else if (instruction_d[6:0] == 7'b1100011 && (
            (instruction_d[14:12] == 3'b000 && zero_flag_e) || // BEQ
            (instruction_d[14:12] == 3'b001 && !zero_flag_e)   // BNE
        )) begin
            // Branch
            pc_next = pc_reg + immediate;
        end else if (instruction_d[6:0] == 7'b1100111) begin
            // JALR
            pc_next = rs1_data_d + immediate;
        end else begin
            // Próxima instrução sequencial
            pc_next = pc_reg + 32'h00000004;
        end
    end
    
    // Interface de memória
    assign mem_data_out = rs2_data_e;
    assign mem_req = mem_we_e || (instruction_f[6:0] == 7'b0000011); // WE ou LW
    
    // PCIe interface
    assign pcie_tx_data = writeback_data_w;
    assign pcie_tx_valid = (wb_sel_m == 2'b10); // Após JAL/JALR
    
    // Saídas de status multiplexadas
    assign status_sel = 4'b0000; // PC value by default
    assign status_data = pc_reg; // Valor fixo para exemplo
    
    // Instância da NPU Top
    npu_top #(
        .DATA_WIDTH(32),
        .ADDR_WIDTH(32)
    ) npu_inst (
        .clk(clk),
        .rst_n(rst_n),
        .bus_addr(mem_addr),
        .bus_data_in(mem_data_in),
        .bus_cmd({mem_we, mem_re, 1'b0}), // Codificação dos comandos
        .bus_ready(mem_ready),
        .bus_data_out(mem_data_out),
        .bus_req(mem_req),
        .mem_addr(),
        .mem_data_out(),
        .mem_we(),
        .mem_re(),
        .mem_data_in(),
        .mem_mem_ready(),
        .ready(),
        .done()
    );

endmodule